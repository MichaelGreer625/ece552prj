module alu
(
    input [15:0] a,
    input [15:0] b,
    input [3:0] control,
    output [15:0] result,
    output [2:0] flags
);



endmodule
