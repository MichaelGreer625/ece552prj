/*
  mode table
  1 0 | OP
  ----------
  0 0 | SLL 
  0 1 | SRA
  1 0 | ROR
  1 1 | *
*/

module shifter
(
    input [15:0] shift_in,
    input [3:0] shift_val
    input [1:0] mode,
    output [15:0] shift_out 
);



endmodule
