module addsub16
(
    input [] a,
    input [] b,
    input sub,
    output [15:0] sum
);



endmodule
